module InstBuffer(
    input wire clk,
    input wire rst
);

endmodule // InstBuffer