`include "defines.v"

module regfile(input wire clk,
               input wire rst,
               input wire we,                  // write or not
               input wire[`RegAddrBus] waddr,
               input wire[`RegBus] wdata,
               input wire re1,                 // write or not
               input wire[`RegAddrBus] raddr1,
               output reg[`RegBus] rdata1,
               input wire re2,                 // write or not
               input wire[`RegAddrBus] raddr2,
               output reg[`RegBus] rdata2);
    
    reg[`RegBus] regs[0:`RegNum-1];
    initial begin
        regs[0] <= `ZeroWord;
        regs[1] <= `ZeroWord;
        regs[2] <= `ZeroWord;
        regs[3] <= `ZeroWord;
        regs[4] <= `ZeroWord;
        regs[5] <= `ZeroWord;
        regs[6] <= `ZeroWord;
        regs[7] <= `ZeroWord;
        regs[8] <= `ZeroWord;
        regs[9] <= `ZeroWord;
        regs[10] <= `ZeroWord;
        regs[11] <= `ZeroWord;
        regs[12] <= `ZeroWord;
        regs[13] <= `ZeroWord;
        regs[14] <= `ZeroWord;
        regs[15] <= `ZeroWord;
        regs[16] <= `ZeroWord;
        regs[17] <= `ZeroWord;
        regs[18] <= `ZeroWord;
        regs[19] <= `ZeroWord;
        regs[20] <= `ZeroWord;
        regs[21] <= `ZeroWord;
        regs[22] <= `ZeroWord;
        regs[23] <= `ZeroWord;
        regs[24] <= `ZeroWord;
        regs[25] <= `ZeroWord;
        regs[26] <= `ZeroWord;
        regs[27] <= `ZeroWord;
        regs[28] <= `ZeroWord;
        regs[29] <= `ZeroWord;
        regs[30] <= `ZeroWord;
        regs[31] <= `ZeroWord;
    end
    
    // genvar i;
    // generate
    // for (i = 0; i < 32; i = i + 1) begin : label
    //     NOTE: Argument inside can only be muodule
    //     instanation
    // end
    // endgenerate
    
    
    // ----------- wirte operation --------------
    always @(posedge clk) begin
        if (rst == `RstDisable) begin
            $display("Answer is ", regs[1]);
            if ((we == `WriteEnable) && (waddr != `RegNumLog2'h0))
            begin
                regs[waddr] <= wdata;
            end
        end
    end
    // ------------ read operation ---------------
    always @(*) begin
        if (rst == `RstEnable || raddr2 == `RegNumLog2'h0) begin
            // Knowing that register 0 is always ZEROWORD
            rdata1 <= `ZeroWord;
            end else if ((raddr1 == waddr) && (we == `WriteEnable) &&
            (re1 == `ReadEnable)) begin
            rdata1 <= wdata;
            end else if (re1 == `ReadEnable) begin
            rdata1 <= regs[raddr1];
            end else begin
            rdata1 <= `ZeroWord;
        end
    end
    
    always @(*) begin
        if (rst == `RstEnable || raddr2 == `RegNumLog2'h0) begin
            rdata2 <= `ZeroWord;
            end else if ((raddr2 == waddr) && (we == `WriteEnable) &&
            (re2 == `ReadEnable)) begin
            rdata2 <= wdata;
            end else if (re2 == `ReadEnable) begin
            rdata2 <= regs[raddr2];
            end else begin
            rdata2 <= `ZeroWord;
        end
    end
    
endmodule // regfile
