// connect to 4 stage module to control stalls
// Possible Improvement 
// 1. out-of-order execution (renaming...)
// 2. multiple issueing (multiple modules to decode )
// 3. data forwarding 
// 4. Cache memory


module StallControler(
    input wire rst,
    input wire clk,
    output wire [31:0] stall
);

endmodule // StallControler